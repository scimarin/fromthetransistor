module control_unit(
    input wire clk, reset,
    output reg write
);
endmodule
