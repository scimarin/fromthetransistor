module cpu_casing();

// links CPU to MMU
// links MMU to TLB
// latches the memory bus

endmodule
