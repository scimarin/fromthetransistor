module computer;
// will contain cpu.v and memory.v
endmodule
