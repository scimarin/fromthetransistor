module computer();

// links the cpu_casing to memory

endmodule
