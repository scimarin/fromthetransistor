module processing_unit();

// contains registers, the bus and the ALU

endmodule
