module cpu(
    input wire clk,
    input wire reset,
    input wire [31:0] from_memory,
    output wire [31:0] address,
    output wire [31:0] to_memory,
    output reg write
);

    data_path _dp(

    );

    control_unit _cu(

    );

endmodule
