module cpu;
endmodule;
