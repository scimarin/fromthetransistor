module memory;
// will contain modules for program ROM memory, data RW memory + stuff from the IO ports
endmodule;
