module shift_register()
